// This file holds the hazard detection unit.

module hazard_unit(
    input 
    output hazard
);

endmodule

