// This file holds the hazard detection unit.

module hazard_unit(
    input clk,
    output hazard
);

endmodule

